module ALU_control(
    ins,
    ALUOp,
    ALUCtrl
);

input  [5:0] ins;
input  [1:0] ALUOp;
output [3:0] ALUCtrl;

endmodule
